.title KiCad schematic
.include "LM4040_NA2P048_TRANS.lib"
RR3 Net-_R3-Pad1_ Net-_Q1-Pad3_ 75
QQ1 Net-_Q1-Pad1_ Net-_Q1-Pad2_ Net-_Q1-Pad3_ 2N7002
UU1 ? Net-_R3-Pad1_ Net-_R5-Pad1_ Net-_R8-Pad1_ NO2 ? VDD Net-_U1-Pad10_ VDD Net-_U1-Pad10_ MICS-4514
RR8 Net-_R8-Pad1_ Net-_Q2-Pad3_ 50
QQ2 Net-_Q2-Pad1_ Net-_Q2-Pad2_ Net-_Q2-Pad3_ 2N7002
CC3 vin GND 22u
RR12 NO2 GNDD 1M
RR11 NO2 Net-_Q6-Pad3_ 100K
PP1 PWM SCALE_1 SCALE_2 CO NO2 CONN_01X05
PP2 GND GNDD VREF VDD vin CONN_01X05
QQ6 SCALE_1 GNDD Net-_Q6-Pad3_ 2N7002
QQ5 SCALE_2 GNDD Net-_Q5-Pad3_ 2N7002
RR9 NO2 Net-_Q5-Pad3_ 10K
RR6 CO GNDD 1M
RR5 Net-_R5-Pad1_ Net-_Q4-Pad3_ 100K
QQ4 SCALE_1 GNDD Net-_Q4-Pad3_ 2N7002
QQ3 SCALE_2 GNDD Net-_Q3-Pad3_ 2N7002
RR4 CO Net-_Q3-Pad3_ 10K
RR7 vin VREF 560
DD1 VREF GNDD LM4040
CC1 VDD GNDD 22u
RR14 VDD vin 100
RR15 GNDD GND 100
RR13 Net-_Q2-Pad2_ GND R
RR2 Net-_Q1-Pad2_ GND R
RR10 PWM Net-_Q2-Pad1_ 47k
RR1 PWM Net-_Q1-Pad1_ 47k
QQ7 Net-_Q1-Pad2_ GND Net-_Q1-Pad1_ BC849
QQ8 Net-_Q2-Pad2_ GND Net-_Q2-Pad1_ BC849
.end
